----------------------------------------------------------------------
-- Project		:	Invent a Chip
-- Authors		:	Jan D�rre
-- Year  		:	2013
-- Description	:	This example tests every 7-seg-display by using 
--					address a counter to generate every possible
--					output. For the 4 hex-displays the counter runs
--					from 0 to 15, for the dec-displays the counter
--					runs from -1000 to 1000. 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.iac_pkg.all;

entity invent_a_chip is
	port (
		-- Global Signals
		clock				: in  std_ulogic;
		reset				: in  std_ulogic;
		-- Interface Signals
		-- 7-Seg
		sevenseg_cs   		: out std_ulogic;
		sevenseg_wr   		: out std_ulogic;
		sevenseg_addr 		: out std_ulogic_vector(CW_ADDR_SEVENSEG-1 downto 0);
		sevenseg_din  		: in  std_ulogic_vector(CW_DATA_SEVENSEG-1 downto 0);
		sevenseg_dout 		: out std_ulogic_vector(CW_DATA_SEVENSEG-1 downto 0);
		-- ADC/DAC
		adc_dac_cs 	 		: out std_ulogic;
		adc_dac_wr 	 		: out std_ulogic;
		adc_dac_addr 		: out std_ulogic_vector(CW_ADDR_ADC_DAC-1 downto 0);
		adc_dac_din  		: in  std_ulogic_vector(CW_DATA_ADC_DAC-1 downto 0);
		adc_dac_dout 		: out std_ulogic_vector(CW_DATA_ADC_DAC-1 downto 0);
		-- AUDIO
		audio_cs   			: out std_ulogic;
		audio_wr   			: out std_ulogic;
		audio_addr 			: out std_ulogic_vector(CW_ADDR_AUDIO-1 downto 0);
		audio_din  			: in  std_ulogic_vector(CW_DATA_AUDIO-1 downto 0);
		audio_dout 			: out std_ulogic_vector(CW_DATA_AUDIO-1 downto 0);
		audio_irq_left  	: in  std_ulogic;
		audio_irq_right 	: in  std_ulogic;
		audio_ack_left  	: out std_ulogic;
		audio_ack_right 	: out std_ulogic;
		-- Infra-red Receiver
		ir_cs				: out std_ulogic;
		ir_wr				: out std_ulogic;
		ir_addr				: out std_ulogic_vector(CW_ADDR_IR-1 downto 0);
		ir_din				: in  std_ulogic_vector(CW_DATA_IR-1 downto 0);
		ir_dout				: out std_ulogic_vector(CW_DATA_IR-1 downto 0);
		ir_irq_rx			: in  std_ulogic;
		ir_ack_rx			: out std_ulogic;
		-- LCD
		lcd_cs   			: out std_ulogic;
		lcd_wr   			: out std_ulogic;
		lcd_addr 			: out std_ulogic_vector(CW_ADDR_LCD-1 downto 0);
		lcd_din  			: in  std_ulogic_vector(CW_DATA_LCD-1 downto 0);
		lcd_dout 			: out std_ulogic_vector(CW_DATA_LCD-1 downto 0);
		lcd_irq_rdy			: in  std_ulogic;
		lcd_ack_rdy			: out std_ulogic;
		-- SRAM
		sram_cs   			: out std_ulogic;
		sram_wr   			: out std_ulogic;
		sram_addr 			: out std_ulogic_vector(CW_ADDR_SRAM-1 downto 0);
		sram_din  			: in  std_ulogic_vector(CW_DATA_SRAM-1 downto 0);
		sram_dout 			: out std_ulogic_vector(CW_DATA_SRAM-1 downto 0);
		-- UART
		uart_cs   	  		: out std_ulogic;
		uart_wr   	  		: out std_ulogic;
		uart_addr 	  		: out std_ulogic_vector(CW_ADDR_UART-1 downto 0);
		uart_din  	  		: in  std_ulogic_vector(CW_DATA_UART-1 downto 0);
		uart_dout 	  		: out std_ulogic_vector(CW_DATA_UART-1 downto 0);
		uart_irq_rx  		: in  std_ulogic;
		uart_irq_tx  		: in  std_ulogic;
		uart_ack_rx  		: out std_ulogic;
		uart_ack_tx  		: out std_ulogic;
		-- GPIO
		gp_ctrl 			: out std_ulogic_vector(15 downto 0);
		gp_in 				: in  std_ulogic_vector(15 downto 0);
		gp_out				: out std_ulogic_vector(15 downto 0);
		-- LED/Switches/Keys
		led_green			: out std_ulogic_vector(8  downto 0);
		led_red				: out std_ulogic_vector(17 downto 0);
		switch				: in  std_ulogic_vector(17 downto 0);
		key 				: in  std_ulogic_vector(2  downto 0)
	);
end invent_a_chip;

architecture rtl of invent_a_chip is

	-- speed
	constant SPEED_RATE : natural := CV_SYS_CLOCK_RATE/16;

	-- state register
	type state_t is (HEX_TEST, DEC_TEST, DO_NOTHING);
	signal state, state_nxt : state_t;
	
	-- counter register for every possible dec-value
	signal cnt, cnt_nxt 			: signed(to_log2(2001)-1 downto 0); -- -1000..0..1000
	
	-- counter for enable signal (SYS_CLOCK/16)
	signal cnt_enable, cnt_enable_nxt 	: unsigned(to_log2(SPEED_RATE)-1 downto 0);
	
	-- enable signal, generated by cnt_enable
	signal enable : std_ulogic;
	
	-- mask for hex displays
	signal hex_mask, hex_mask_nxt : std_ulogic_vector(3 downto 0);

begin

	-- sequential process
	process (clock, reset)
	begin
		-- async reset
		if reset = '1' then
			state 		<= HEX_TEST;
			cnt 		<= (others => '0');
			cnt_enable	<= (others => '0');
			hex_mask 	<= "0001";
		elsif rising_edge(clock) then	
			state 		<= state_nxt;
			cnt 		<= cnt_nxt;
			cnt_enable	<= cnt_enable_nxt;
			hex_mask 	<= hex_mask_nxt;
		end if;
	end process;
	
	
	-- logic for enable generator
	process (cnt_enable)
	begin
		if cnt_enable >= to_unsigned(SPEED_RATE, cnt_enable'length) then
			cnt_enable_nxt 	<= (others => '0');
			enable 			<= '1';
		else
			cnt_enable_nxt <= cnt_enable + to_unsigned(1, cnt_enable'length);
			enable 			<= '0';
		end if;
	end process;
	
	
	-- logic
	process (state, cnt, enable, hex_mask)
	begin
		-- standard assignments
		
		-- hold values of registers
		state_nxt 	  	<= state;
		cnt_nxt 	  	<= cnt;
		hex_mask_nxt 	<= hex_mask;
		
		-- set bus signals to standard values (not in use)
		sevenseg_cs		<= '0';
		sevenseg_wr		<= '0';
		sevenseg_addr	<= (others => '0');
		sevenseg_dout	<= (others => '0');
		
		
		-- turn of leds
		led_green	<= (others => '0');
		led_red		<= (others => '0');
		
		-- state machine
		case state is
			-- starting state
			when HEX_TEST =>
				-- indicate state HEX_TEST
				led_green(0) <= '1';
				
				-- for every possible hex-value
				if cnt <= to_signed(15, cnt'length) then
					
					-- wait for enable signal
					if enable = '1' then
						-- set chip select for seven-segment-interface
						sevenseg_cs <= '1';
						-- set write mode
						sevenseg_wr <= '1';
						-- set address, use mask to select hex-display, LSB has to be zero for hexmode
						sevenseg_addr <= std_ulogic_vector(resize(unsigned(hex_mask & '0'), sevenseg_addr'length));
						-- set data (4 times cnt-value)
						sevenseg_dout <= std_ulogic_vector(resize(unsigned(cnt(3 downto 0) & cnt(3 downto 0) & cnt(3 downto 0) & cnt(3 downto 0)), sevenseg_dout'length));
						
						-- inc counter
						cnt_nxt <= cnt + to_signed(1, cnt'length);
					end if;
					
				else
				
					-- last mask not reached
					if hex_mask(3) = '0' then
					
						-- shift mask
						hex_mask_nxt <= std_ulogic_vector(shift_left(unsigned(hex_mask), 1));
						
						-- reset counter
						cnt_nxt <= (others => '0');
					
					else
						-- next state
						state_nxt <= DEC_TEST;
				
						-- reset counter
						cnt_nxt <= to_signed(-1000, cnt'length);
					end if;
				
				end if;
				
			-- test every value from -1000 to 1000 (-1000 and 1000 should produce error on display)
			when DEC_TEST => 
				-- indicate state DEC_TEST
				led_green(1) <= '1';
				
				-- wait for enable signal
				if enable = '1' then
					-- set chip select for seven-segment-interface
					sevenseg_cs <= '1';
					-- set write mode
					sevenseg_wr <= '1';
					-- set address
					sevenseg_addr <= CV_ADDR_SEVENSEG_DEC;
					-- set data
					sevenseg_dout <= std_ulogic_vector(resize(cnt, sevenseg_dout'length));
					
					-- end cnt reached
					if cnt = to_signed(1000, cnt'length) then 
						-- end test
						state_nxt <= DO_NOTHING;
					else
						-- inc counter
						cnt_nxt <= signed(cnt) + to_signed(1, cnt'length);
					end if;
				end if;
			
			-- wait forever
			when DO_NOTHING =>
				-- indicate state DO_NOTHING
				led_green(2) <= '1';
			
		end case;
	end process;
	
	-- default assignments for unused signals
	gp_ctrl 			<= (others => '0');
	gp_out				<= (others => '0');	
	adc_dac_cs 	 		<= '0';
	adc_dac_wr 	 		<= '0';
	adc_dac_addr 		<= (others => '0');
	adc_dac_dout 		<= (others => '0');
	audio_cs 	 		<= '0';
	audio_wr 	 		<= '0';
	audio_addr 	 		<= (others => '0');
	audio_dout 	 		<= (others => '0');
	audio_ack_left  	<= '0';
	audio_ack_right 	<= '0';
	ir_cs				<= '0';
	ir_wr				<= '0';
	ir_addr				<= (others => '0');
	ir_dout				<= (others => '0');
	ir_ack_rx			<= '0';
	lcd_cs 	 	 		<= '0';
	lcd_wr 	 	 		<= '0';
	lcd_addr 	 		<= (others => '0');
	lcd_dout 	 		<= (others => '0');
	lcd_ack_rdy			<= '0';
	sram_cs 	 		<= '0';
	sram_wr 	 		<= '0';
	sram_addr 	 		<= (others => '0');
	sram_dout 	 		<= (others => '0');
	uart_cs 	 		<= '0';
	uart_wr 	 		<= '0';
	uart_addr 	 		<= (others => '0');
	uart_dout 	 		<= (others => '0');
	uart_ack_rx  		<= '0';
	uart_ack_tx  		<= '0';

end rtl;